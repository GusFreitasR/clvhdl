library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library KAILIB;

package regBank_states is
    
	TYPE Regbank_states IS (IDLE, pickingReg, reading, writing);

	 
end package regBank_states;